/*
 *
 */

module datapath (
	input         coreclk   ,
	input         core_arstn,
	dfi_if.master m_dfi
);

	

endmodule // datapath
