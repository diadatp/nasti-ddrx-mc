
typedef enum logic [1:0] {c9 = 2'b00, c10, c11} col_widths;
typedef enum logic [2:0] {r11 = 3'b000, r12, r13, r14, r15} row_widths;
