

`define C_NASTI_ID_WIDTH   9
`define C_NASTI_ADDR_WIDTH 32
`define C_NASTI_DATA_WIDTH 64
`define C_NASTI_USER_WIDTH 1
`define C_NASTILITE_ADDR_WIDTH 6
`define C_NASTILITE_DATA_WIDTH 64
