/**
 *
 */

module nastilite_frontend (
    input              s_nastilite_clk    ,
    input              s_nastilite_aresetn,
    nastilite_if.slave s_nastilite
);

endmodule