/*
 *
 */

module phy_top (
    // DDR PHY Interface
    input         dfi_clk    ,
    input         dfi_clkdiv2,
    input         dfi_clkdiv4,
    input         dfi_arstn  ,
    dfi_if.slave  s_dfi      ,
    // DDR3 Interface
    inout  [63:0] ddr_dq     ,
    output [ 7:0] ddr_dqs_n  ,
    output [ 7:0] ddr_dqs_p  ,
    output [15:0] ddr_addr   ,
    output [ 2:0] ddr_ba     ,
    output        ddr_ras_n  ,
    output        ddr_cas_n  ,
    output        ddr_we_n   ,
    output        ddr_reset_n,
    output [ 1:0] ddr_ck_p   ,
    output [ 1:0] ddr_ck_n   ,
    output [ 1:0] ddr_cke    ,
    output [ 1:0] ddr_cs_n   ,
    output [ 7:0] ddr_dm     ,
    output [ 1:0] ddr_odt
);

    logic dfi_arst = ~dfi_arstn;

    OBUFT #(
        .DRIVE     (12       ), // Specify the output drive strength
        .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
        .SLEW      ("SLOW"   )  // Specify the output slew rate
    ) ras_n_OBUFT_inst (
        .O(ddr_ras_n      ), // Buffer output (connect directly to top-level port)
        .I(s_dfi.dfi_ras_n), // Buffer input
        .T(1'b0           )  // 3-state enable input
    );

    OBUFT #(
        .DRIVE     (12       ), // Specify the output drive strength
        .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
        .SLEW      ("SLOW"   )  // Specify the output slew rate
    ) cas_n_OBUFT_inst (
        .O(ddr_cas_n      ), // Buffer output (connect directly to top-level port)
        .I(s_dfi.dfi_cas_n), // Buffer input
        .T(1'b0           )  // 3-state enable input
    );

    OBUFT #(
        .DRIVE     (12       ), // Specify the output drive strength
        .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
        .SLEW      ("SLOW"   )  // Specify the output slew rate
    ) reset_n_OBUFT_inst (
        .O(ddr_reset_n      ), // Buffer output (connect directly to top-level port)
        .I(s_dfi.dfi_reset_n), // Buffer input
        .T(1'b0             )  // 3-state enable input
    );

    OBUFT #(
        .DRIVE     (12       ), // Specify the output drive strength
        .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
        .SLEW      ("SLOW"   )  // Specify the output slew rate
    ) we_n_OBUFT_inst (
        .O(ddr_we_n      ), // Buffer output (connect directly to top-level port)
        .I(s_dfi.dfi_we_n), // Buffer input
        .T(1'b0          )  // 3-state enable input
    );

    generate
        for (genvar ba_i = 0; ba_i < 3; ba_i++) begin : gen_ba
            OBUFT #(
                .DRIVE     (12       ), // Specify the output drive strength
                .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
                .SLEW      ("SLOW"   )  // Specify the output slew rate
            ) ba_OBUFT_inst (
                .O(ddr_ba[ba_i]        ), // Buffer output (connect directly to top-level port)
                .I(s_dfi.dfi_bank[ba_i]), // Buffer input
                .T(1'b0                )  // 3-state enable input
            );
        end
    endgenerate

    generate
        for (genvar addr_i = 0; addr_i < 16; addr_i++) begin : gen_addr
            OBUFT #(
                .DRIVE     (12       ), // Specify the output drive strength
                .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
                .SLEW      ("SLOW"   )  // Specify the output slew rate
            ) addr_OBUFT_inst (
                .O(ddr_addr[addr_i]         ), // Buffer output (connect directly to top-level port)
                .I(s_dfi.dfi_address[addr_i]), // Buffer input
                .T(1'b0                     )  // 3-state enable input
            );
        end
    endgenerate

    generate
        for (genvar cke_i = 0; cke_i < 2; cke_i++) begin : gen_cke
            OBUFT #(
                .DRIVE     (12       ), // Specify the output drive strength
                .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
                .SLEW      ("SLOW"   )  // Specify the output slew rate
            ) cke_OBUFT_inst (
                .O(ddr_cke[cke_i]      ), // Buffer output (connect directly to top-level port)
                .I(s_dfi.dfi_cke[cke_i]), // Buffer input
                .T(1'b0                )  // 3-state enable input
            );
        end
    endgenerate

    generate
        for (genvar cs_n_i = 0; cs_n_i < 2; cs_n_i++) begin : gen_cs_n
            OBUFT #(
                .DRIVE     (12       ), // Specify the output drive strength
                .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
                .SLEW      ("SLOW"   )  // Specify the output slew rate
            ) _OBUFT_inst (
                .O(ddr_cs_n[cs_n_i]      ), // Buffer output (connect directly to top-level port)
                .I(s_dfi.dfi_cs_n[cs_n_i]), // Buffer input
                .T(1'b0                  )  // 3-state enable input
            );
        end
    endgenerate

    generate
        for (genvar dm_i = 0; dm_i < 8; dm_i++) begin : gen_dm
            OBUFT #(
                .DRIVE     (12       ), // Specify the output drive strength
                .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
                .SLEW      ("SLOW"   )  // Specify the output slew rate
            ) dm_OBUFT_inst (
                .O(ddr_dm[dm_i]               ), // Buffer output (connect directly to top-level port)
                .I(s_dfi.dfi_wrdata_mask[dm_i]), // Buffer input
                .T(1'b0                       )  // 3-state enable input
            );
        end
    endgenerate

    generate
        for (genvar odt_i = 0; odt_i < 2; odt_i++) begin : gen_odt
            OBUFT #(
                .DRIVE     (12       ), // Specify the output drive strength
                .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
                .SLEW      ("SLOW"   )  // Specify the output slew rate
            ) odt_OBUFT_inst (
                .O(ddr_odt[odt_i]      ), // Buffer output (connect directly to top-level port)
                .I(s_dfi.dfi_odt[odt_i]), // Buffer input
                .T(1'b0                )  // 3-state enable input
            );
        end
    endgenerate

    logic dq_oser_rst;

    logic [7:0][7:0] dq_odly_cntout;
    logic [7:0][7:0] dq_odly_ce    ;
    logic [7:0][7:0] dq_odly_cntin ;
    logic [7:0][7:0] dq_odly_ld    ;
    logic [7:0][7:0] dq_odly_inc   ;

    logic [7:0][7:0] dq_idly_cntout;
    logic [7:0][7:0] dq_idly_ce    ;
    logic [7:0][7:0] dq_idly_cntin ;
    logic [7:0][7:0] dq_idly_ld    ;
    logic [7:0][7:0] dq_idly_inc   ;

    logic dq_iobuf_dci;
    logic dq_iobuf_id ;
    logic dq_iobuf_t  ;

    logic [7:0] out_fifo_aempty;
    logic [7:0] out_fifo_afull ;
    logic [7:0] out_fifo_empty ;
    logic [7:0] out_fifo_full  ;
    logic       out_fifo_rden  ;

    generate
        for (genvar io_fifo_i = 0; io_fifo_i < 8; io_fifo_i++) begin : gen_io_fifo

            logic [7:0][3:0] out_fifo_q;
            logic [7:0][7:0] out_fifo_d;

            logic [7:0][3:0] dq_iser_q;
            logic [7:0][7:0] in_fifo_q;

            OUT_FIFO #(
                .ALMOST_EMPTY_VALUE(1                 ), // Almost empty offset (1-2)
                .ALMOST_FULL_VALUE (1                 ), // Almost full offset (1-2)
                .ARRAY_MODE        ("ARRAY_MODE_8_X_4"), // ARRAY_MODE_8_X_4, ARRAY_MODE_4_X_4
                .OUTPUT_DISABLE    ("FALSE"           ), // Disable output (FALSE, TRUE)
                .SYNCHRONOUS_MODE  ("FALSE"           )  // Must always be set to false.
            ) OUT_FIFO_inst (
                // FIFO Status Flags: 1-bit (each) output: Flags and other FIFO status outputs
                .ALMOSTEMPTY(out_fifo_aempty[io_fifo_i]), // 1-bit output: Almost empty flag
                .ALMOSTFULL (out_fifo_afull[io_fifo_i] ), // 1-bit output: Almost full flag
                .EMPTY      (out_fifo_empty[io_fifo_i] ), // 1-bit output: Empty flag
                .FULL       (out_fifo_full[io_fifo_i]  ), // 1-bit output: Full flag
                // Q0-Q9: 4-bit (each) output: FIFO Outputs
                .Q0         (out_fifo_q[0]             ), // 4-bit output: Channel 0 output bus
                .Q1         (out_fifo_q[1]             ), // 4-bit output: Channel 1 output bus
                .Q2         (out_fifo_q[2]             ), // 4-bit output: Channel 2 output bus
                .Q3         (out_fifo_q[3]             ), // 4-bit output: Channel 3 output bus
                .Q4         (out_fifo_q[4]             ), // 4-bit output: Channel 4 output bus
                .Q5         (out_fifo_q[5]             ), // 8-bit output: Channel 5 output bus
                .Q6         (out_fifo_q[6]             ), // 8-bit output: Channel 6 output bus
                .Q7         (out_fifo_q[7]             ), // 4-bit output: Channel 7 output bus
                .Q8         (                          ), // 4-bit output: Channel 8 output bus
                .Q9         (                          ), // 4-bit output: Channel 9 output bus
                // D0-D9: 8-bit (each) input: FIFO inputs
                .D0         (out_fifo_d[0]             ), // 8-bit input: Channel 0 input bus
                .D1         (out_fifo_d[1]             ), // 8-bit input: Channel 1 input bus
                .D2         (out_fifo_d[2]             ), // 8-bit input: Channel 2 input bus
                .D3         (out_fifo_d[3]             ), // 8-bit input: Channel 3 input bus
                .D4         (out_fifo_d[4]             ), // 8-bit input: Channel 4 input bus
                .D5         (out_fifo_d[5]             ), // 8-bit input: Channel 5 input bus
                .D6         (out_fifo_d[6]             ), // 8-bit input: Channel 6 input bus
                .D7         (out_fifo_d[7]             ), // 8-bit input: Channel 7 input bus
                .D8         (                          ), // 8-bit input: Channel 8 input bus
                .D9         (                          ), // 8-bit input: Channel 9 input bus
                // FIFO Control Signals: 1-bit (each) input: Clocks, Resets and Enables
                .RDCLK      (dfi_clkdiv4               ), // 1-bit input: Read clock
                .RDEN       (out_fifo_rden             ), // 1-bit input: Read enable
                .RESET      (out_fifo_reset            ), // 1-bit input: Active high reset
                .WRCLK      (                          ), // 1-bit input: Write clock
                .WREN       (                          )  // 1-bit input: Write enable
            );

            IN_FIFO #(
                .ALMOST_EMPTY_VALUE(1                 ), // Almost empty offset (1-2)
                .ALMOST_FULL_VALUE (1                 ), // Almost full offset (1-2)
                .ARRAY_MODE        ("ARRAY_MODE_4_X_8"), // ARRAY_MODE_4_X_8, ARRAY_MODE_4_X_4
                .SYNCHRONOUS_MODE  ("FALSE"           )  // Clock synchronous (FALSE)
            ) IN_FIFO_inst (
                // FIFO Status Flags: 1-bit (each) output: Flags and other FIFO status outputs
                .ALMOSTEMPTY(            ), // 1-bit output: Almost empty
                .ALMOSTFULL (            ), // 1-bit output: Almost full
                .EMPTY      (            ), // 1-bit output: Empty
                .FULL       (            ), // 1-bit output: Full
                // Q0-Q9: 8-bit (each) output: FIFO Outputs
                .Q0         (in_fifo_q[0]), // 8-bit output: Channel 0
                .Q1         (in_fifo_q[1]), // 8-bit output: Channel 1
                .Q2         (in_fifo_q[2]), // 8-bit output: Channel 2
                .Q3         (in_fifo_q[3]), // 8-bit output: Channel 3
                .Q4         (in_fifo_q[4]), // 8-bit output: Channel 4
                .Q5         (in_fifo_q[5]), // 8-bit output: Channel 5
                .Q6         (in_fifo_q[6]), // 8-bit output: Channel 6
                .Q7         (in_fifo_q[7]), // 8-bit output: Channel 7
                .Q8         (            ), // 8-bit output: Channel 8
                .Q9         (            ), // 8-bit output: Channel 9
                // D0-D9: 4-bit (each) input: FIFO inputs
                .D0         (dq_iser_q[0]), // 4-bit input: Channel 0
                .D1         (dq_iser_q[1]), // 4-bit input: Channel 1
                .D2         (dq_iser_q[2]), // 4-bit input: Channel 2
                .D3         (dq_iser_q[3]), // 4-bit input: Channel 3
                .D4         (dq_iser_q[4]), // 4-bit input: Channel 4
                .D5         (dq_iser_q[5]), // 8-bit input: Channel 5
                .D6         (dq_iser_q[6]), // 8-bit input: Channel 6
                .D7         (dq_iser_q[7]), // 4-bit input: Channel 7
                .D8         (            ), // 4-bit input: Channel 8
                .D9         (            ), // 4-bit input: Channel 9
                // FIFO Control Signals: 1-bit (each) input: Clocks, Resets and Enables
                .RDCLK      (            ), // 1-bit input: Read clock
                .RDEN       (            ), // 1-bit input: Read enable
                .RESET      (in_fifo_rst ), // 1-bit input: Reset
                .WRCLK      (            ), // 1-bit input: Write clock
                .WREN       (            )  // 1-bit input: Write enable
            );

            for (genvar dq_i = 0; dq_i < 8; dq_i++) begin : gen_dq

                logic dq_oser_ofb;
                logic dq_in      ;
                logic dq_delayed ;

                OSERDESE2 #(
                    .DATA_RATE_OQ  ("DDR"   ), // DDR, SDR
                    .DATA_RATE_TQ  ("DDR"   ), // DDR, BUF, SDR
                    .DATA_WIDTH    (4       ), // Parallel data width (2-8,10,14)
                    .INIT_OQ       (1'b0    ), // Initial value of OQ output (1'b0,1'b1)
                    .INIT_TQ       (1'b0    ), // Initial value of TQ output (1'b0,1'b1)
                    .SERDES_MODE   ("MASTER"), // MASTER, SLAVE
                    .SRVAL_OQ      (1'b0    ), // OQ output value when SR is used (1'b0,1'b1)
                    .SRVAL_TQ      (1'b0    ), // TQ output value when SR is used (1'b0,1'b1)
                    .TBYTE_CTL     ("FALSE" ), // Enable tristate byte operation (FALSE, TRUE)
                    .TBYTE_SRC     ("FALSE" ), // Tristate byte source (FALSE, TRUE)
                    .TRISTATE_WIDTH(4       )  // 3-state converter width (1,4)
                ) OSERDESE2_inst (
                    .OFB      (dq_oser_ofb          ), // 1-bit output: Feedback path for data
                    .OQ       (                     ), // 1-bit output: Data path output
                    // SHIFTOUT1 / SHIFTOUT2: 1-bit (each) output: Data output expansion (1-bit each)
                    .SHIFTOUT1(                     ),
                    .SHIFTOUT2(                     ),
                    .TBYTEOUT (                     ), // 1-bit output: Byte group tristate
                    .TFB      (                     ), // 1-bit output: 3-state control
                    .TQ       (                     ), // 1-bit output: 3-state control
                    .CLK      (dfi_clk              ), // 1-bit input: High speed clock
                    .CLKDIV   (dfi_clkdiv2          ), // 1-bit input: Divided clock
                    // D1 - D8: 1-bit (each) input: Parallel data inputs (1-bit each)
                    .D1       (out_fifo_q[dq_i%8][0]),
                    .D2       (out_fifo_q[dq_i%8][1]),
                    .D3       (out_fifo_q[dq_i%8][2]),
                    .D4       (out_fifo_q[dq_i%8][3]),
                    .D5       (                     ),
                    .D6       (                     ),
                    .D7       (                     ),
                    .D8       (                     ),
                    .OCE      (1'b1                 ), // 1-bit input: Output data clock enable
                    .RST      (dq_oser_rst          ), // 1-bit input: Reset
                    // SHIFTIN1 / SHIFTIN2: 1-bit (each) input: Data input expansion (1-bit each)
                    .SHIFTIN1 (                     ),
                    .SHIFTIN2 (                     ),
                    // T1 - T4: 1-bit (each) input: Parallel 3-state inputs
                    .T1       (                     ),
                    .T2       (                     ),
                    .T3       (                     ),
                    .T4       (                     ),
                    .TBYTEIN  (                     ), // 1-bit input: Byte group tristate
                    .TCE      (                     )  // 1-bit input: 3-state clock enable
                );

                (* IODELAY_GROUP = "dq_iodelay_group" *) // Specifies group name for associated IDELAYs/ODELAYs and IDELAYCTRL

                    ODELAYE2 #(
                        .CINVCTRL_SEL         ("FALSE"   ), // Enable dynamic clock inversion (FALSE, TRUE)
                        .DELAY_SRC            ("ODATAIN" ), // Delay input (ODATAIN, CLKIN)
                        .HIGH_PERFORMANCE_MODE("TRUE"    ), // Reduced jitter ("TRUE"), Reduced power ("FALSE")
                        .ODELAY_TYPE          ("VAR_LOAD"), // FIXED, VARIABLE, VAR_LOAD, VAR_LOAD_PIPE
                        .ODELAY_VALUE         (0         ), // Output delay tap setting (0-31)
                        .PIPE_SEL             ("FALSE"   ), // Select pipelined mode, FALSE, TRUE
                        .REFCLK_FREQUENCY     (200.0     ), // IDELAYCTRL clock input frequency in MHz (190.0-210.0, 290.0-310.0).
                        .SIGNAL_PATTERN       ("DATA"    )  // DATA, CLOCK input signal
                    ) ODELAYE2_inst (
                        .CNTVALUEOUT(dq_odly_cntout[io_fifo_i][dq_i]), // 5-bit output: Counter value output
                        .DATAOUT    (dq_delayed                     ), // 1-bit output: Delayed data/clock output
                        .C          (dfi_clkdiv4                    ), // 1-bit input: Clock input
                        .CE         (dq_odly_ce[io_fifo_i][dq_i]    ), // 1-bit input: Active high enable increment/decrement input
                        .CINVCTRL   (1'b0                           ), // 1-bit input: Dynamic clock inversion input
                        .CLKIN      (1'b0                           ), // 1-bit input: Clock delay input
                        .CNTVALUEIN (dq_odly_cntin[io_fifo_i][dq_i] ), // 5-bit input: Counter value input
                        .INC        (dq_odly_inc[io_fifo_i][dq_i]   ), // 1-bit input: Increment / Decrement tap delay input
                        .LD         (dq_odly_ld[io_fifo_i][dq_i]    ), // 1-bit input: Loads ODELAY_VALUE tap delay in VARIABLE mode, in VAR_LOAD or VAR_LOAD_PIPE mode, loads the value of CNTVALUEIN
                        .LDPIPEEN   (1'b0                           ), // 1-bit input: Enables the pipeline register to load data
                        .ODATAIN    (dq_oser_ofb                    ), // 1-bit input: Output delay data input
                        .REGRST     (dq_odly_rst                    )  // 1-bit input: Active-high reset tap-delay input
                    );

                ISERDESE2 #(
                    .DATA_RATE        ("DDR"   ), // DDR, SDR
                    .DATA_WIDTH       (4       ), // Parallel data width (2-8,10,14)
                    .DYN_CLKDIV_INV_EN("FALSE" ), // Enable DYNCLKDIVINVSEL inversion (FALSE, TRUE)
                    .DYN_CLK_INV_EN   ("FALSE" ), // Enable DYNCLKINVSEL inversion (FALSE, TRUE)
                    // INIT_Q1 - INIT_Q4: Initial value on the Q outputs (0/1)
                    .INIT_Q1          (1'b0    ),
                    .INIT_Q2          (1'b0    ),
                    .INIT_Q3          (1'b0    ),
                    .INIT_Q4          (1'b0    ),
                    .INTERFACE_TYPE   ("MEMORY"), // MEMORY, MEMORY_DDR3, MEMORY_QDR, NETWORKING, OVERSAMPLE
                    .IOBDELAY         ("BOTH"  ), // NONE, BOTH, IBUF, IFD
                    .NUM_CE           (2       ), // Number of clock enables (1,2)
                    .OFB_USED         ("FALSE" ), // Select OFB path (FALSE, TRUE)
                    .SERDES_MODE      ("MASTER"), // MASTER, SLAVE
                    // SRVAL_Q1 - SRVAL_Q4: Q output values when SR is used (0/1)
                    .SRVAL_Q1         (1'b0    ),
                    .SRVAL_Q2         (1'b0    ),
                    .SRVAL_Q3         (1'b0    ),
                    .SRVAL_Q4         (1'b0    )
                ) ISERDESE2_inst (
                    .O           (                      ), // 1-bit output: Combinatorial output
                    // Q1 - Q8: 1-bit (each) output: Registered data outputs
                    .Q1          (dq_iser_q[dq_i%8][0]  ),
                    .Q2          (dq_iser_q[dq_i%8][1]  ),
                    .Q3          (dq_iser_q[dq_i%8][2]  ),
                    .Q4          (dq_iser_q[dq_i%8][3]  ),
                    .Q5          (                      ),
                    .Q6          (                      ),
                    .Q7          (                      ),
                    .Q8          (                      ),
                    // SHIFTOUT1, SHIFTOUT2: 1-bit (each) output: Data width expansion output ports
                    .SHIFTOUT1   (                      ),
                    .SHIFTOUT2   (                      ),
                    .BITSLIP     (1'b0                  ), // 1-bit input: The BITSLIP pin performs a Bitslip operation synchronous to
                    // CLKDIV when asserted (active High). Subsequently, the data seen on the Q1
                    // to Q8 output ports will shift, as in a barrel-shifter operation, one
                    // position every time Bitslip is invoked (DDR operation is different from
                    // SDR).
                    
                    // CE1, CE2: 1-bit (each) input: Data register clock enable inputs
                    .CE1         (1'b1                  ),
                    .CE2         (1'b1                  ),
                    .CLKDIVP     (                      ), // 1-bit input: TBD
                    // Clocks: 1-bit (each) input: ISERDESE2 clock input ports
                    .CLK         (dqs_bufio_p[in_fifo_i]), // 1-bit input: High-speed clock
                    .CLKB        (dqs_bufio_n[in_fifo_i]), // 1-bit input: High-speed secondary clock
                    .CLKDIV      (dfi_clkdiv2           ), // 1-bit input: Divided clock
                    .OCLK        (dfi_clk               ), // 1-bit input: High speed output clock used when INTERFACE_TYPE="MEMORY"
                    // Dynamic Clock Inversions: 1-bit (each) input: Dynamic clock inversion pins to switch clock polarity
                    .DYNCLKDIVSEL(                      ), // 1-bit input: Dynamic CLKDIV inversion
                    .DYNCLKSEL   (                      ), // 1-bit input: Dynamic CLK/CLKB inversion
                    // Input Data: 1-bit (each) input: ISERDESE2 data input ports
                    .D           (1'b0                  ), // 1-bit input: Data input
                    .DDLY        (dq_in_delayed         ), // 1-bit input: Serial data from IDELAYE2
                    .OFB         (                      ), // 1-bit input: Data feedback from OSERDESE2
                    .OCLKB       (                      ), // 1-bit input: High speed negative edge output clock
                    .RST         (dq_iser_rst           ), // 1-bit input: Active high asynchronous reset
                    // SHIFTIN1, SHIFTIN2: 1-bit (each) input: Data width expansion input ports
                    .SHIFTIN1    (                      ),
                    .SHIFTIN2    (                      )
                );

                (* IODELAY_GROUP = "dq_iodelay_group" *) // Specifies group name for associated IDELAYs/ODELAYs and IDELAYCTRL

                    IDELAYE2 #(
                        .CINVCTRL_SEL         ("FALSE"   ), // Enable dynamic clock inversion (FALSE, TRUE)
                        .DELAY_SRC            ("IDATAIN" ), // Delay input (IDATAIN, DATAIN)
                        .HIGH_PERFORMANCE_MODE("TRUE"    ), // Reduced jitter ("TRUE"), Reduced power ("FALSE")
                        .IDELAY_TYPE          ("VAR_LOAD"), // FIXED, VARIABLE, VAR_LOAD, VAR_LOAD_PIPE
                        .IDELAY_VALUE         (0         ), // Input delay tap setting (0-31)
                        .PIPE_SEL             ("FALSE"   ), // Select pipelined mode, FALSE, TRUE
                        .REFCLK_FREQUENCY     (200.0     ), // IDELAYCTRL clock input frequency in MHz (190.0-210.0, 290.0-310.0).
                        .SIGNAL_PATTERN       ("DATA"    )  // DATA, CLOCK input signal
                    ) IDELAYE2_inst (
                        .CNTVALUEOUT(dq_idly_cntout[io_fifo_i][dq_i]), // 5-bit output: Counter value output
                        .DATAOUT    (dq_in_delayed                  ), // 1-bit output: Delayed data output
                        .C          (dfi_clkdiv4                    ), // 1-bit input: Clock input
                        .CE         (dq_idly_ce[io_fifo_i][dq_i]    ), // 1-bit input: Active high enable increment/decrement input
                        .CINVCTRL   (1'b0                           ), // 1-bit input: Dynamic clock inversion input
                        .CNTVALUEIN (dq_idly_cntin[io_fifo_i][dq_i] ), // 5-bit input: Counter value input
                        .DATAIN     (1'b0                           ), // 1-bit input: Internal delay data input
                        .IDATAIN    (dq_in                          ), // 1-bit input: Data input from the I/O
                        .INC        (dq_idly_inc[io_fifo_i][dq_i]   ), // 1-bit input: Increment / Decrement tap delay input
                        .LD         (dq_idly_ld[io_fifo_i][dq_i]    ), // 1-bit input: Load IDELAY_VALUE input
                        .LDPIPEEN   (1'b0                           ), // 1-bit input: Enable PIPELINE register to load data input
                        .REGRST     (dq_idly_rst                    )  // 1-bit input: Active-high reset tap-delay input
                    );

                IOBUF_DCIEN #(
                    .DRIVE          (12            ), // Specify the output drive strength
                    .IBUF_LOW_PWR   ("TRUE"        ), // Low Power - "TRUE", High Performance = "FALSE"
                    .IOSTANDARD     ("SSTL15_T_DCI"), // Specify the I/O standard
                    .SLEW           ("SLOW"        ), // Specify the output slew rate
                    .USE_IBUFDISABLE("TRUE"        )  // Use IBUFDISABLE function, "TRUE" or "FALSE"
                ) IOBUF_DCIEN_inst (
                    .O             (dq_in       ), // Buffer output
                    .IO            (ddr_dq[dq_i]), // Buffer inout port (connect directly to top-level port)
                    .DCITERMDISABLE(dq_iobuf_dci), // DCI Termination enable input
                    .I             (dq_delayed  ), // Buffer input
                    .IBUFDISABLE   (dq_iobuf_id ), // Input disable input, low=disable
                    .T             (dq_iobuf_t  )  // 3-state enable input, high=input, low=output
                );

            end
        end
    endgenerate

    logic dqs_oddr_rst;

    logic [7:0] dqs_bufio_p;
    logic [7:0] dqs_bufio_n;

    logic [7:0] dqs_iobuf_tm ;
    logic [7:0] dqs_iobuf_ts ;
    logic [7:0] dqs_iobuf_dci;
    logic [7:0] dqs_iobuf_id ;
    logic [7:0] dqs_iobuf_t  ;

    logic [7:0] dqs_idly_cntout;
    logic [7:0] dqs_idly_ce    ;
    logic [7:0] dqs_idly_cntin ;
    logic [7:0] dqs_idly_ld    ;
    logic [7:0] dqs_idly_inc   ;

    logic [7:0] dqs_odly_cntout;
    logic [7:0] dqs_odly_ce    ;
    logic [7:0] dqs_odly_cntin ;
    logic [7:0] dqs_odly_ld    ;
    logic [7:0] dqs_odly_inc   ;

    (* IODELAY_GROUP = "dqs_iodelay_group" *) // Specifies group name for associated IDELAYs/ODELAYs and IDELAYCTRL

        IDELAYCTRL IDELAYCTRL_inst (
            .RDY   (dqs_idlyctrl_rdy), // 1-bit output: Ready output
            .REFCLK(dfi_clkdiv4     ), // 1-bit input: Reference clock input
            .RST   (dqs_idlyctrl_rst)  // 1-bit input: Active high reset input
        );

    generate
        for (genvar dqs_i = 0; dqs_i < 8; dqs_i++) begin : gen_dqs

            logic dqs_oddr        ;
            logic dqs_in_delayed_p;
            logic dqs_in_delayed_n;
            logic dqs_in_p        ;
            logic dqs_in_n        ;

            ODDR #(
                .DDR_CLK_EDGE("SAME_EDGE"), // "OPPOSITE_EDGE" or "SAME_EDGE"
                .INIT        (1'b0       ), // Initial value of Q: 1'b0 or 1'b1
                .SRTYPE      ("SYNC"     )  // Set/Reset type: "SYNC" or "ASYNC"
            ) ODDR_inst (
                .Q (dqs_oddr    ), // 1-bit DDR output
                .C (dfi_clk     ), // 1-bit clock input
                .CE(1'b1        ), // 1-bit clock enable input
                .D1(1'b1        ), // 1-bit data input (positive edge)
                .D2(1'b0        ), // 1-bit data input (negative edge)
                .R (dqs_oddr_rst), // 1-bit reset
                .S (1'b0        )  // 1-bit set
            );

            (* IODELAY_GROUP = "dqs_iodelay_group" *) // Specifies group name for associated IDELAYs/ODELAYs and IDELAYCTRL

                IDELAYE2 #(
                    .CINVCTRL_SEL         ("FALSE"   ), // Enable dynamic clock inversion (FALSE, TRUE)
                    .DELAY_SRC            ("IDATAIN" ), // Delay input (IDATAIN, DATAIN)
                    .HIGH_PERFORMANCE_MODE("TRUE"    ), // Reduced jitter ("TRUE"), Reduced power ("FALSE")
                    .IDELAY_TYPE          ("VAR_LOAD"), // FIXED, VARIABLE, VAR_LOAD, VAR_LOAD_PIPE
                    .IDELAY_VALUE         (0         ), // Input delay tap setting (0-31)
                    .PIPE_SEL             ("FALSE"   ), // Select pipelined mode, FALSE, TRUE
                    .REFCLK_FREQUENCY     (200.0     ), // IDELAYCTRL clock input frequency in MHz (190.0-210.0, 290.0-310.0).
                    .SIGNAL_PATTERN       ("DATA"    )  // DATA, CLOCK input signal
                ) IDELAYE2_inst_p (
                    .CNTVALUEOUT(dqs_idly_cntout[dqs_i]), // 5-bit output: Counter value output
                    .DATAOUT    (dqs_in_delayed_p      ), // 1-bit output: Delayed data output
                    .C          (dfi_clkdiv4           ), // 1-bit input: Clock input
                    .CE         (dqs_idly_ce[dqs_i]    ), // 1-bit input: Active high enable increment/decrement input
                    .CINVCTRL   (1'b0                  ), // 1-bit input: Dynamic clock inversion input
                    .CNTVALUEIN (dqs_idly_cntin[dqs_i] ), // 5-bit input: Counter value input
                    .DATAIN     (1'b0                  ), // 1-bit input: Internal delay data input
                    .IDATAIN    (dqs_in_p              ), // 1-bit input: Data input from the I/O
                    .INC        (dqs_idly_inc[dqs_i]   ), // 1-bit input: Increment / Decrement tap delay input
                    .LD         (dqs_idly_ld[dqs_i]    ), // 1-bit input: Load IDELAY_VALUE input
                    .LDPIPEEN   (1'b0                  ), // 1-bit input: Enable PIPELINE register to load data input
                    .REGRST     (dqs_idly_rst          )  // 1-bit input: Active-high reset tap-delay input
                );

            (* IODELAY_GROUP = "dqs_iodelay_group" *) // Specifies group name for associated IDELAYs/ODELAYs and IDELAYCTRL

                IDELAYE2 #(
                    .CINVCTRL_SEL         ("FALSE"   ), // Enable dynamic clock inversion (FALSE, TRUE)
                    .DELAY_SRC            ("IDATAIN" ), // Delay input (IDATAIN, DATAIN)
                    .HIGH_PERFORMANCE_MODE("TRUE"    ), // Reduced jitter ("TRUE"), Reduced power ("FALSE")
                    .IDELAY_TYPE          ("VAR_LOAD"), // FIXED, VARIABLE, VAR_LOAD, VAR_LOAD_PIPE
                    .IDELAY_VALUE         (0         ), // Input delay tap setting (0-31)
                    .PIPE_SEL             ("FALSE"   ), // Select pipelined mode, FALSE, TRUE
                    .REFCLK_FREQUENCY     (200.0     ), // IDELAYCTRL clock input frequency in MHz (190.0-210.0, 290.0-310.0).
                    .SIGNAL_PATTERN       ("DATA"    )  // DATA, CLOCK input signal
                ) IDELAYE2_inst_n (
                    .CNTVALUEOUT(dqs_idly_cntout[dqs_i]), // 5-bit output: Counter value output
                    .DATAOUT    (dqs_in_delayed_n        ), // 1-bit output: Delayed data output
                    .C          (dfi_clkdiv4           ), // 1-bit input: Clock input
                    .CE         (dqs_idly_ce[dqs_i]    ), // 1-bit input: Active high enable increment/decrement input
                    .CINVCTRL   (1'b0                  ), // 1-bit input: Dynamic clock inversion input
                    .CNTVALUEIN (dqs_idly_cntin[dqs_i] ), // 5-bit input: Counter value input
                    .DATAIN     (1'b0                  ), // 1-bit input: Internal delay data input
                    .IDATAIN    (dqs_in_n              ), // 1-bit input: Data input from the I/O
                    .INC        (dqs_idly_inc[dqs_i]   ), // 1-bit input: Increment / Decrement tap delay input
                    .LD         (dqs_idly_ld[dqs_i]    ), // 1-bit input: Load IDELAY_VALUE input
                    .LDPIPEEN   (1'b0                  ), // 1-bit input: Enable PIPELINE register to load data input
                    .REGRST     (dqs_idly_rst          )  // 1-bit input: Active-high reset tap-delay input
                );

            BUFIO BUFIO_inst_p (
                .O(dqs_bufio_p[dqs_i]), // 1-bit output: Clock output (connect to I/O clock loads).
                .I(dqs_in_delayed_p  )  // 1-bit input: Clock input (connect to an IBUFG or BUFMR).
            );

            BUFIO BUFIO_inst_n (
                .O(dqs_bufio_n[dqs_i]), // 1-bit output: Clock output (connect to I/O clock loads).
                .I(dqs_in_delayed_n  )  // 1-bit input: Clock input (connect to an IBUFG or BUFMR).
            );

            (* IODELAY_GROUP = "dqs_iodelay_group" *) // Specifies group name for associated IDELAYs/ODELAYs and IDELAYCTRL

                ODELAYE2 #(
                    .CINVCTRL_SEL         ("FALSE"   ), // Enable dynamic clock inversion (FALSE, TRUE)
                    .DELAY_SRC            ("ODATAIN" ), // Delay input (ODATAIN, CLKIN)
                    .HIGH_PERFORMANCE_MODE("TRUE"    ), // Reduced jitter ("TRUE"), Reduced power ("FALSE")
                    .ODELAY_TYPE          ("VAR_LOAD"), // FIXED, VARIABLE, VAR_LOAD, VAR_LOAD_PIPE
                    .ODELAY_VALUE         (0         ), // Output delay tap setting (0-31)
                    .PIPE_SEL             ("FALSE"   ), // Select pipelined mode, FALSE, TRUE
                    .REFCLK_FREQUENCY     (200.0     ), // IDELAYCTRL clock input frequency in MHz (190.0-210.0, 290.0-310.0).
                    .SIGNAL_PATTERN       ("DATA"    )  // DATA, CLOCK input signal
                ) ODELAYE2_inst (
                    .CNTVALUEOUT(dqs_odly_cntout[dqs_i]), // 5-bit output: Counter value output
                    .DATAOUT    (dqs_delayed           ), // 1-bit output: Delayed data/clock output
                    .C          (dfi_clkdiv4           ), // 1-bit input: Clock input
                    .CE         (dqs_odly_ce[dqs_i]    ), // 1-bit input: Active high enable increment/decrement input
                    .CINVCTRL   (1'b0                  ), // 1-bit input: Dynamic clock inversion input
                    .CLKIN      (1'b0                  ), // 1-bit input: Clock delay input
                    .CNTVALUEIN (dqs_odly_cntin[dqs_i] ), // 5-bit input: Counter value input
                    .INC        (dqs_odly_inc[dqs_i]   ), // 1-bit input: Increment / Decrement tap delay input
                    .LD         (dqs_odly_ld[dqs_i]    ), // 1-bit input: Loads ODELAY_VALUE tap delay in VARIABLE mode, in VAR_LOAD or VAR_LOAD_PIPE mode, loads the value of CNTVALUEIN
                    .LDPIPEEN   (1'b0                  ), // 1-bit input: Enables the pipeline register to load data
                    .ODATAIN    (dqs_oddr              ), // 1-bit input: Output delay data input
                    .REGRST     (dqs_odly_rst          )  // 1-bit input: Active-high reset tap-delay input
                );

            IOBUFDS_DIFF_OUT_DCIEN #(
                .DIFF_TERM      ("FALSE"            ), // Differential Termination ("TRUE"/"FALSE")
                .IBUF_LOW_PWR   ("FALSE"            ), // Low Power - "TRUE", High Performance = "FALSE"
                .IOSTANDARD     ("DIFF_SSTL15_T_DCI"), // Specify the I/O standard
                .USE_IBUFDISABLE("TRUE"             )  // Use IBUFDISABLE function, "TRUE" or "FALSE"
            ) IOBUFDS_DIFF_OUT_DCIEN_inst (
                .O             (dqs_in_p            ), // Buffer p-side output
                .OB            (dqs_in_n            ), // Buffer n-side output
                .IO            (ddr_dqs_p[dqs_i]    ), // Diff_p inout (connect directly to top-level port)
                .IOB           (ddr_dqs_n[dqs_i]    ), // Diff_n inout (connect directly to top-level port)
                .DCITERMDISABLE(dqs_iobuf_dci[dqs_i]), // DCI Termination enable input
                .I             (dqs_delayed         ), // Buffer input
                .IBUFDISABLE   (dqs_iobuf_id[dqs_i] ), // Input disable input, high=disable
                .TM            (dqs_iobuf_tm[dqs_i] ), // 3-state enable input, high=input, low=output
                .TS            (dqs_iobuf_ts[dqs_i] )  // 3-state enable input, high=input, low=output
            );

        end
    endgenerate

    generate
        for (genvar ddr_ck_i = 0; ddr_ck_i < 2; ddr_ck_i++) begin : gen_ck

            logic ddr_ck;

            ODDR #(
                .DDR_CLK_EDGE("SAME_EDGE"), // "OPPOSITE_EDGE" or "SAME_EDGE"
                .INIT        (1'b0       ), // Initial value of Q: 1'b0 or 1'b1
                .SRTYPE      ("ASYNC"    )  // Set/Reset type: "SYNC" or "ASYNC"
            ) ODDR_inst (
                .Q (ddr_ck  ), // 1-bit DDR output
                .C (dfi_clk ), // 1-bit clock input
                .CE(1'b1    ), // 1-bit clock enable input
                .D1(1'b1    ), // 1-bit data input (positive edge)
                .D2(1'b0    ), // 1-bit data input (negative edge)
                .R (dfi_arst), // 1-bit reset
                .S (1'b0    )  // 1-bit set
            );

            OBUFTDS #(
                .IOSTANDARD("DEFAULT"), // Specify the output I/O standard
                .SLEW      ("SLOW"   )  // Specify the output slew rate
            ) OBUFTDS_inst (
                .O (ddr_ck_p[ddr_ck_i]), // Diff_p output (connect directly to top-level port)
                .OB(ddr_ck_n[ddr_ck_i]), // Diff_n output (connect directly to top-level port)
                .I (ddr_ck            ), // Buffer input
                .T (1'b0              )  // 3-state enable input
            );

        end
    endgenerate

endmodule // phy_top
