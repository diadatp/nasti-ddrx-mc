/*
 *
 */

module datapath (
	input coreclk   ,
	input core_arstn
);

endmodule // datapath
